
`ifndef TEMPLATE_SVH
`define TEMPLATE_SVH


`include "template_transfer.sv"
`include "template_config.sv"

`include "template_master_driver.svh"
`include "template_master_monitor.svh"
`include "template_master_sequencer.svh"
`include "template_master_agent.svh"

`include "template_slave_driver.svh"
`include "template_slave_monitor.svh"
`include "template_slave_sequencer.svh"
`include "template_slave_agent.svh"


`include "template_master_driver.sv"       
`include "template_master_monitor.sv"
`include "template_master_sequencer.sv"
`include "template_master_agent.sv"
`include "template_master_seq_lib.sv"

`include "template_slave_driver.sv"       
`include "template_slave_monitor.sv"
`include "template_slave_sequencer.sv"
`include "template_slave_agent.sv"
`include "template_slave_seq_lib.sv"



   
`endif //  `ifndef TEMPLATE_SVH
