
`ifndef TEMPLATE_SLAVE_SEQUENCER_SV
`define TEMPLATE_SLAVE_SEQUENCER_SV

function template_slave_sequencer::new (string name, uvm_component parent);
  super.new(name, parent);
endfunction : new

`endif // TEMPLATE_SLAVE_SEQUENCER_SV


